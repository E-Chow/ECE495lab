entity bsr_unit is
port(clk, left_right: in std_logic; 
	right_in, left_in: in std_logic;
	q: out std_logic);
end bsr_unit;
